// This is the unpowered netlist.
module tiny_user_project (user_clock2,
    wb_clk_i,
    wb_rst_i,
    wbs_ack_o,
    wbs_cyc_i,
    wbs_stb_i,
    wbs_we_i,
    io_in,
    io_oeb,
    io_out,
    la_data_in,
    la_data_out,
    la_oenb,
    user_irq,
    wbs_adr_i,
    wbs_dat_i,
    wbs_dat_o,
    wbs_sel_i);
 input user_clock2;
 input wb_clk_i;
 input wb_rst_i;
 output wbs_ack_o;
 input wbs_cyc_i;
 input wbs_stb_i;
 input wbs_we_i;
 input [37:0] io_in;
 output [37:0] io_oeb;
 output [37:0] io_out;
 input [63:0] la_data_in;
 output [63:0] la_data_out;
 input [63:0] la_oenb;
 output [2:0] user_irq;
 input [31:0] wbs_adr_i;
 input [31:0] wbs_dat_i;
 output [31:0] wbs_dat_o;
 input [3:0] wbs_sel_i;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire net14;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net15;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net16;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net52;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net53;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net54;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net86;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net87;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net88;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net89;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net90;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net91;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net155;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net156;
 wire net184;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;

 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _019_ (.A1(net4),
    .A2(net3),
    .Z(_000_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _020_ (.A1(net6),
    .A2(net5),
    .A3(_000_),
    .Z(_001_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _021_ (.A1(net1),
    .A2(net2),
    .Z(_002_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _022_ (.A1(net8),
    .A2(net7),
    .A3(_002_),
    .Z(_003_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _023_ (.A1(_001_),
    .A2(_003_),
    .ZN(_004_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _024_ (.A1(net4),
    .A2(net3),
    .B1(net6),
    .B2(net5),
    .ZN(_005_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _025_ (.A1(net4),
    .A2(net3),
    .B1(net6),
    .B2(net5),
    .ZN(_006_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _026_ (.A1(net4),
    .A2(net3),
    .A3(net6),
    .A4(net5),
    .Z(_007_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _027_ (.A1(_005_),
    .A2(_006_),
    .B(_007_),
    .ZN(_008_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _028_ (.A1(net1),
    .A2(net2),
    .B1(net8),
    .B2(net7),
    .ZN(_009_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _029_ (.A1(net1),
    .A2(net2),
    .B1(net8),
    .B2(net7),
    .ZN(_010_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _030_ (.A1(net1),
    .A2(net2),
    .A3(net8),
    .A4(net7),
    .Z(_011_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _031_ (.A1(_009_),
    .A2(_010_),
    .B(_011_),
    .ZN(_012_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _032_ (.A1(_008_),
    .A2(_012_),
    .ZN(_013_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _033_ (.A1(_004_),
    .A2(_013_),
    .Z(_014_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _034_ (.I(_014_),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _035_ (.A1(_007_),
    .A2(_011_),
    .Z(_015_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _036_ (.I(_015_),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _037_ (.A1(_007_),
    .A2(_011_),
    .ZN(_016_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _038_ (.A1(_008_),
    .A2(_012_),
    .ZN(_017_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _039_ (.A1(_004_),
    .A2(_013_),
    .B1(net12),
    .B2(_016_),
    .C(_017_),
    .ZN(net11));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _040_ (.A1(_001_),
    .A2(_003_),
    .Z(_018_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _041_ (.I(_018_),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_14 (.ZN(net14));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_15 (.ZN(net15));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_16 (.ZN(net16));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_17 (.ZN(net17));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_18 (.ZN(net18));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_19 (.ZN(net19));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_20 (.ZN(net20));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_21 (.ZN(net21));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_22 (.ZN(net22));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_23 (.ZN(net23));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_24 (.ZN(net24));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_25 (.ZN(net25));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_26 (.ZN(net26));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_27 (.ZN(net27));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_28 (.ZN(net28));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_29 (.ZN(net29));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_30 (.ZN(net30));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_31 (.ZN(net31));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_32 (.ZN(net32));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_33 (.ZN(net33));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_34 (.ZN(net34));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_35 (.ZN(net35));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_36 (.ZN(net36));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_37 (.ZN(net37));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_38 (.ZN(net38));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_39 (.ZN(net39));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_40 (.ZN(net40));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_41 (.ZN(net41));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_42 (.ZN(net42));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_43 (.ZN(net43));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_44 (.ZN(net44));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_45 (.ZN(net45));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_46 (.ZN(net46));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_47 (.ZN(net47));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_48 (.ZN(net48));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_49 (.ZN(net49));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_50 (.ZN(net50));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_51 (.ZN(net51));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_52 (.ZN(net52));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_53 (.ZN(net53));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_54 (.ZN(net54));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_55 (.ZN(net55));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_56 (.ZN(net56));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_57 (.ZN(net57));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_58 (.ZN(net58));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_59 (.ZN(net59));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_60 (.ZN(net60));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_61 (.ZN(net61));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_62 (.ZN(net62));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_63 (.ZN(net63));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_64 (.ZN(net64));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_65 (.ZN(net65));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_66 (.ZN(net66));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_67 (.ZN(net67));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_68 (.ZN(net68));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_69 (.ZN(net69));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_70 (.ZN(net70));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_71 (.ZN(net71));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_72 (.ZN(net72));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_73 (.ZN(net73));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_74 (.ZN(net74));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_75 (.ZN(net75));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_76 (.ZN(net76));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_77 (.ZN(net77));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_78 (.ZN(net78));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_79 (.ZN(net79));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_80 (.ZN(net80));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_81 (.ZN(net81));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_82 (.ZN(net82));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_83 (.ZN(net83));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_84 (.ZN(net84));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_85 (.ZN(net85));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_86 (.ZN(net86));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_87 (.ZN(net87));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_88 (.ZN(net88));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_89 (.ZN(net89));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_90 (.ZN(net90));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_91 (.ZN(net91));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_92 (.ZN(net92));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_93 (.ZN(net93));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_94 (.ZN(net94));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_95 (.ZN(net95));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_96 (.ZN(net96));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_97 (.ZN(net97));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_98 (.ZN(net98));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_99 (.ZN(net99));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_100 (.ZN(net100));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_101 (.ZN(net101));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_102 (.ZN(net102));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_103 (.ZN(net103));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_104 (.ZN(net104));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_105 (.ZN(net105));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_106 (.ZN(net106));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_107 (.ZN(net107));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_108 (.ZN(net108));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_109 (.ZN(net109));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_110 (.ZN(net110));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_111 (.ZN(net111));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_112 (.ZN(net112));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_113 (.ZN(net113));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_114 (.ZN(net114));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_115 (.ZN(net115));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_116 (.ZN(net116));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_117 (.ZN(net117));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_118 (.ZN(net118));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_119 (.ZN(net119));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_120 (.ZN(net120));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_121 (.ZN(net121));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_122 (.ZN(net122));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_123 (.ZN(net123));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_124 (.ZN(net124));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_125 (.ZN(net125));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_126 (.ZN(net126));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_127 (.ZN(net127));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_128 (.ZN(net128));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_129 (.ZN(net129));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_130 (.ZN(net130));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_131 (.ZN(net131));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_132 (.ZN(net132));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_133 (.ZN(net133));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_134 (.ZN(net134));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_135 (.ZN(net135));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_136 (.ZN(net136));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_137 (.ZN(net137));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_138 (.ZN(net138));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_139 (.ZN(net139));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_140 (.ZN(net140));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_141 (.ZN(net141));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_142 (.ZN(net142));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_143 (.ZN(net143));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_144 (.ZN(net144));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_145 (.ZN(net145));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_146 (.ZN(net146));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_147 (.ZN(net147));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_148 (.ZN(net148));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_149 (.ZN(net149));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_150 (.ZN(net150));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_151 (.ZN(net151));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_152 (.ZN(net152));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_153 (.ZN(net153));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_154 (.ZN(net154));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_155 (.ZN(net155));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_156 (.ZN(net156));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_157 (.ZN(net157));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_158 (.ZN(net158));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_159 (.ZN(net159));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_160 (.ZN(net160));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_161 (.ZN(net161));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_162 (.ZN(net162));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_163 (.ZN(net163));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_164 (.ZN(net164));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_165 (.ZN(net165));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_166 (.ZN(net166));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_167 (.ZN(net167));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_168 (.ZN(net168));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_169 (.ZN(net169));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_170 (.ZN(net170));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_171 (.ZN(net171));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_172 (.ZN(net172));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_173 (.ZN(net173));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_174 (.ZN(net174));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_175 (.ZN(net175));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_176 (.ZN(net176));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_177 (.ZN(net177));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_178 (.ZN(net178));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_179 (.ZN(net179));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_180 (.ZN(net180));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_181 (.ZN(net181));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_182 (.ZN(net182));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_183 (.ZN(net183));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_184 (.ZN(net184));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__037__A1 (.I(_007_));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_9 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_136 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_137 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_138 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_139 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_140 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_141 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_142 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_143 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_144 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_145 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_146 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_147 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_148 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_149 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_150 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_151 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_152 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_153 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_154 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_155 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_156 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_157 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_158 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_159 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_160 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_161 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_162 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_163 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_164 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_165 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_166 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_167 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_168 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_169 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_170 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_171 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_172 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_173 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_174 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_175 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_176 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_177 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_178 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_179 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_180 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_181 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_182 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_183 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_184 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_185 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_186 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_187 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_188 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_189 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_190 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_191 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_192 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_193 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_194 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_195 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_196 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_197 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_198 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_199 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_200 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_201 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_202 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_203 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_204 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_205 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_206 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_207 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_208 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_209 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_210 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_211 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_212 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_213 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_214 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_215 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_216 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_217 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_218 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_219 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_220 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_221 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_222 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_223 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_224 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_225 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_226 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_227 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_228 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_229 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_230 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_231 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_232 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_233 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_234 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_235 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_236 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_237 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_238 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_239 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_240 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_241 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_242 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_243 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_244 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_245 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_246 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_247 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_248 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_249 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_250 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_251 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_252 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_253 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_254 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_255 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_256 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_257 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_258 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_259 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_260 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_261 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_262 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_263 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_264 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_265 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_266 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_267 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_268 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_269 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_270 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_271 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_272 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_273 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_274 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_275 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_276 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_277 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_278 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_279 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_280 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_281 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_282 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_283 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_284 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_285 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_286 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_287 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_288 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_289 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_290 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_291 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_292 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_293 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_294 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_295 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_296 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_297 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_298 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_299 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_300 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_301 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_302 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_303 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_304 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_305 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_306 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_307 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_308 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_309 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_310 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_311 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_312 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_313 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_314 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_315 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_316 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_317 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_318 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_319 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_320 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_321 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_322 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_323 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_324 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_325 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_326 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_327 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_328 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2750 ();
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1 (.I(io_in[10]),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input2 (.I(io_in[11]),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input3 (.I(io_in[12]),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input4 (.I(io_in[13]),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input5 (.I(io_in[14]),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input6 (.I(io_in[15]),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_1 input7 (.I(io_in[8]),
    .Z(net7));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_1 input8 (.I(io_in[9]),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output9 (.I(net9),
    .Z(io_out[16]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output10 (.I(net10),
    .Z(io_out[17]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output11 (.I(net11),
    .Z(io_out[18]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output12 (.I(net12),
    .Z(io_out[19]));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_13 (.ZN(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__035__A1 (.I(_007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__027__B (.I(_007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__037__A2 (.I(_011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__035__A2 (.I(_011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__031__B (.I(_011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(io_in[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(io_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input4_I (.I(io_in[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input5_I (.I(io_in[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input6_I (.I(io_in[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input7_I (.I(io_in[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input8_I (.I(io_in[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__030__A1 (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__029__A1 (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__028__A1 (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__021__A1 (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__030__A2 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__029__A2 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__028__A2 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__021__A2 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__026__A2 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__025__A2 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__024__A2 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__019__A2 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__026__A1 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__025__A1 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__024__A1 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__019__A1 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__026__A4 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__025__B2 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__024__B2 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__020__A2 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__026__A3 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__025__B1 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__024__B1 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__020__A1 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__030__A4 (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__029__B2 (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__028__B2 (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__022__A2 (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output9_I (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output10_I (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output11_I (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output12_I (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__039__B1 (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_19_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_23_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_25_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_29_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_33_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_131_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_133_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_137_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_139_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_141_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_145_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_145_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_146_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_146_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_147_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_147_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_148_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_149_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_149_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_150_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_150_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_151_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_151_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_152_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_152_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_153_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_153_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_154_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_154_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_155_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_155_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_156_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_156_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_157_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_157_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_158_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_158_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_158_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_159_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_159_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_160_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_160_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_161_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_161_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_162_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_163_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_163_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_164_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_164_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_164_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_164_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_164_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1043 ();
 assign io_oeb[0] = net13;
 assign io_oeb[10] = net23;
 assign io_oeb[11] = net24;
 assign io_oeb[12] = net25;
 assign io_oeb[13] = net26;
 assign io_oeb[14] = net27;
 assign io_oeb[15] = net28;
 assign io_oeb[16] = net29;
 assign io_oeb[17] = net30;
 assign io_oeb[18] = net31;
 assign io_oeb[19] = net32;
 assign io_oeb[1] = net14;
 assign io_oeb[20] = net33;
 assign io_oeb[21] = net34;
 assign io_oeb[22] = net35;
 assign io_oeb[23] = net36;
 assign io_oeb[24] = net37;
 assign io_oeb[25] = net38;
 assign io_oeb[26] = net39;
 assign io_oeb[27] = net40;
 assign io_oeb[28] = net41;
 assign io_oeb[29] = net42;
 assign io_oeb[2] = net15;
 assign io_oeb[30] = net43;
 assign io_oeb[31] = net44;
 assign io_oeb[32] = net45;
 assign io_oeb[33] = net46;
 assign io_oeb[34] = net47;
 assign io_oeb[35] = net48;
 assign io_oeb[36] = net49;
 assign io_oeb[37] = net50;
 assign io_oeb[3] = net16;
 assign io_oeb[4] = net17;
 assign io_oeb[5] = net18;
 assign io_oeb[6] = net19;
 assign io_oeb[7] = net20;
 assign io_oeb[8] = net21;
 assign io_oeb[9] = net22;
 assign io_out[0] = net51;
 assign io_out[10] = net61;
 assign io_out[11] = net62;
 assign io_out[12] = net63;
 assign io_out[13] = net64;
 assign io_out[14] = net65;
 assign io_out[15] = net66;
 assign io_out[1] = net52;
 assign io_out[20] = net67;
 assign io_out[21] = net68;
 assign io_out[22] = net69;
 assign io_out[23] = net70;
 assign io_out[24] = net71;
 assign io_out[25] = net72;
 assign io_out[26] = net73;
 assign io_out[27] = net74;
 assign io_out[28] = net75;
 assign io_out[29] = net76;
 assign io_out[2] = net53;
 assign io_out[30] = net77;
 assign io_out[31] = net78;
 assign io_out[32] = net79;
 assign io_out[33] = net80;
 assign io_out[34] = net81;
 assign io_out[35] = net82;
 assign io_out[36] = net83;
 assign io_out[37] = net84;
 assign io_out[3] = net54;
 assign io_out[4] = net55;
 assign io_out[5] = net56;
 assign io_out[6] = net57;
 assign io_out[7] = net58;
 assign io_out[8] = net59;
 assign io_out[9] = net60;
 assign la_data_out[0] = net85;
 assign la_data_out[10] = net95;
 assign la_data_out[11] = net96;
 assign la_data_out[12] = net97;
 assign la_data_out[13] = net98;
 assign la_data_out[14] = net99;
 assign la_data_out[15] = net100;
 assign la_data_out[16] = net101;
 assign la_data_out[17] = net102;
 assign la_data_out[18] = net103;
 assign la_data_out[19] = net104;
 assign la_data_out[1] = net86;
 assign la_data_out[20] = net105;
 assign la_data_out[21] = net106;
 assign la_data_out[22] = net107;
 assign la_data_out[23] = net108;
 assign la_data_out[24] = net109;
 assign la_data_out[25] = net110;
 assign la_data_out[26] = net111;
 assign la_data_out[27] = net112;
 assign la_data_out[28] = net113;
 assign la_data_out[29] = net114;
 assign la_data_out[2] = net87;
 assign la_data_out[30] = net115;
 assign la_data_out[31] = net116;
 assign la_data_out[32] = net117;
 assign la_data_out[33] = net118;
 assign la_data_out[34] = net119;
 assign la_data_out[35] = net120;
 assign la_data_out[36] = net121;
 assign la_data_out[37] = net122;
 assign la_data_out[38] = net123;
 assign la_data_out[39] = net124;
 assign la_data_out[3] = net88;
 assign la_data_out[40] = net125;
 assign la_data_out[41] = net126;
 assign la_data_out[42] = net127;
 assign la_data_out[43] = net128;
 assign la_data_out[44] = net129;
 assign la_data_out[45] = net130;
 assign la_data_out[46] = net131;
 assign la_data_out[47] = net132;
 assign la_data_out[48] = net133;
 assign la_data_out[49] = net134;
 assign la_data_out[4] = net89;
 assign la_data_out[50] = net135;
 assign la_data_out[51] = net136;
 assign la_data_out[52] = net137;
 assign la_data_out[53] = net138;
 assign la_data_out[54] = net139;
 assign la_data_out[55] = net140;
 assign la_data_out[56] = net141;
 assign la_data_out[57] = net142;
 assign la_data_out[58] = net143;
 assign la_data_out[59] = net144;
 assign la_data_out[5] = net90;
 assign la_data_out[60] = net145;
 assign la_data_out[61] = net146;
 assign la_data_out[62] = net147;
 assign la_data_out[63] = net148;
 assign la_data_out[6] = net91;
 assign la_data_out[7] = net92;
 assign la_data_out[8] = net93;
 assign la_data_out[9] = net94;
 assign user_irq[0] = net149;
 assign user_irq[1] = net150;
 assign user_irq[2] = net151;
 assign wbs_ack_o = net152;
 assign wbs_dat_o[0] = net153;
 assign wbs_dat_o[10] = net163;
 assign wbs_dat_o[11] = net164;
 assign wbs_dat_o[12] = net165;
 assign wbs_dat_o[13] = net166;
 assign wbs_dat_o[14] = net167;
 assign wbs_dat_o[15] = net168;
 assign wbs_dat_o[16] = net169;
 assign wbs_dat_o[17] = net170;
 assign wbs_dat_o[18] = net171;
 assign wbs_dat_o[19] = net172;
 assign wbs_dat_o[1] = net154;
 assign wbs_dat_o[20] = net173;
 assign wbs_dat_o[21] = net174;
 assign wbs_dat_o[22] = net175;
 assign wbs_dat_o[23] = net176;
 assign wbs_dat_o[24] = net177;
 assign wbs_dat_o[25] = net178;
 assign wbs_dat_o[26] = net179;
 assign wbs_dat_o[27] = net180;
 assign wbs_dat_o[28] = net181;
 assign wbs_dat_o[29] = net182;
 assign wbs_dat_o[2] = net155;
 assign wbs_dat_o[30] = net183;
 assign wbs_dat_o[31] = net184;
 assign wbs_dat_o[3] = net156;
 assign wbs_dat_o[4] = net157;
 assign wbs_dat_o[5] = net158;
 assign wbs_dat_o[6] = net159;
 assign wbs_dat_o[7] = net160;
 assign wbs_dat_o[8] = net161;
 assign wbs_dat_o[9] = net162;
endmodule

