magic
tech gf180mcuC
magscale 1 5
timestamp 1670229143
<< obsm1 >>
rect 672 855 59304 66345
<< metal2 >>
rect 0 67600 56 67900
rect 672 67600 728 67900
rect 1344 67600 1400 67900
rect 2016 67600 2072 67900
rect 2688 67600 2744 67900
rect 3360 67600 3416 67900
rect 3696 67600 3752 67900
rect 4368 67600 4424 67900
rect 5040 67600 5096 67900
rect 5712 67600 5768 67900
rect 6384 67600 6440 67900
rect 7056 67600 7112 67900
rect 7392 67600 7448 67900
rect 8064 67600 8120 67900
rect 8736 67600 8792 67900
rect 9408 67600 9464 67900
rect 10080 67600 10136 67900
rect 10752 67600 10808 67900
rect 11088 67600 11144 67900
rect 11760 67600 11816 67900
rect 12432 67600 12488 67900
rect 13104 67600 13160 67900
rect 13776 67600 13832 67900
rect 14448 67600 14504 67900
rect 14784 67600 14840 67900
rect 15456 67600 15512 67900
rect 16128 67600 16184 67900
rect 16800 67600 16856 67900
rect 17472 67600 17528 67900
rect 18144 67600 18200 67900
rect 18480 67600 18536 67900
rect 19152 67600 19208 67900
rect 19824 67600 19880 67900
rect 20496 67600 20552 67900
rect 21168 67600 21224 67900
rect 21840 67600 21896 67900
rect 22176 67600 22232 67900
rect 22848 67600 22904 67900
rect 23520 67600 23576 67900
rect 24192 67600 24248 67900
rect 24864 67600 24920 67900
rect 25536 67600 25592 67900
rect 25872 67600 25928 67900
rect 26544 67600 26600 67900
rect 27216 67600 27272 67900
rect 27888 67600 27944 67900
rect 28560 67600 28616 67900
rect 29232 67600 29288 67900
rect 29904 67600 29960 67900
rect 30240 67600 30296 67900
rect 30912 67600 30968 67900
rect 31584 67600 31640 67900
rect 32256 67600 32312 67900
rect 32928 67600 32984 67900
rect 33600 67600 33656 67900
rect 33936 67600 33992 67900
rect 34608 67600 34664 67900
rect 35280 67600 35336 67900
rect 35952 67600 36008 67900
rect 36624 67600 36680 67900
rect 37296 67600 37352 67900
rect 37632 67600 37688 67900
rect 38304 67600 38360 67900
rect 38976 67600 39032 67900
rect 39648 67600 39704 67900
rect 40320 67600 40376 67900
rect 40992 67600 41048 67900
rect 41328 67600 41384 67900
rect 42000 67600 42056 67900
rect 42672 67600 42728 67900
rect 43344 67600 43400 67900
rect 44016 67600 44072 67900
rect 44688 67600 44744 67900
rect 45024 67600 45080 67900
rect 45696 67600 45752 67900
rect 46368 67600 46424 67900
rect 47040 67600 47096 67900
rect 47712 67600 47768 67900
rect 48384 67600 48440 67900
rect 48720 67600 48776 67900
rect 49392 67600 49448 67900
rect 50064 67600 50120 67900
rect 50736 67600 50792 67900
rect 51408 67600 51464 67900
rect 52080 67600 52136 67900
rect 52416 67600 52472 67900
rect 53088 67600 53144 67900
rect 53760 67600 53816 67900
rect 54432 67600 54488 67900
rect 55104 67600 55160 67900
rect 55776 67600 55832 67900
rect 56112 67600 56168 67900
rect 56784 67600 56840 67900
rect 57456 67600 57512 67900
rect 58128 67600 58184 67900
rect 58800 67600 58856 67900
rect 59472 67600 59528 67900
rect 59808 67600 59864 67900
rect 0 100 56 400
rect 336 100 392 400
rect 1008 100 1064 400
rect 1680 100 1736 400
rect 2352 100 2408 400
rect 3024 100 3080 400
rect 3696 100 3752 400
rect 4032 100 4088 400
rect 4704 100 4760 400
rect 5376 100 5432 400
rect 6048 100 6104 400
rect 6720 100 6776 400
rect 7392 100 7448 400
rect 7728 100 7784 400
rect 8400 100 8456 400
rect 9072 100 9128 400
rect 9744 100 9800 400
rect 10416 100 10472 400
rect 11088 100 11144 400
rect 11424 100 11480 400
rect 12096 100 12152 400
rect 12768 100 12824 400
rect 13440 100 13496 400
rect 14112 100 14168 400
rect 14784 100 14840 400
rect 15120 100 15176 400
rect 15792 100 15848 400
rect 16464 100 16520 400
rect 17136 100 17192 400
rect 17808 100 17864 400
rect 18480 100 18536 400
rect 18816 100 18872 400
rect 19488 100 19544 400
rect 20160 100 20216 400
rect 20832 100 20888 400
rect 21504 100 21560 400
rect 22176 100 22232 400
rect 22512 100 22568 400
rect 23184 100 23240 400
rect 23856 100 23912 400
rect 24528 100 24584 400
rect 25200 100 25256 400
rect 25872 100 25928 400
rect 26208 100 26264 400
rect 26880 100 26936 400
rect 27552 100 27608 400
rect 28224 100 28280 400
rect 28896 100 28952 400
rect 29568 100 29624 400
rect 29904 100 29960 400
rect 30576 100 30632 400
rect 31248 100 31304 400
rect 31920 100 31976 400
rect 32592 100 32648 400
rect 33264 100 33320 400
rect 33936 100 33992 400
rect 34272 100 34328 400
rect 34944 100 35000 400
rect 35616 100 35672 400
rect 36288 100 36344 400
rect 36960 100 37016 400
rect 37632 100 37688 400
rect 37968 100 38024 400
rect 38640 100 38696 400
rect 39312 100 39368 400
rect 39984 100 40040 400
rect 40656 100 40712 400
rect 41328 100 41384 400
rect 41664 100 41720 400
rect 42336 100 42392 400
rect 43008 100 43064 400
rect 43680 100 43736 400
rect 44352 100 44408 400
rect 45024 100 45080 400
rect 45360 100 45416 400
rect 46032 100 46088 400
rect 46704 100 46760 400
rect 47376 100 47432 400
rect 48048 100 48104 400
rect 48720 100 48776 400
rect 49056 100 49112 400
rect 49728 100 49784 400
rect 50400 100 50456 400
rect 51072 100 51128 400
rect 51744 100 51800 400
rect 52416 100 52472 400
rect 52752 100 52808 400
rect 53424 100 53480 400
rect 54096 100 54152 400
rect 54768 100 54824 400
rect 55440 100 55496 400
rect 56112 100 56168 400
rect 56448 100 56504 400
rect 57120 100 57176 400
rect 57792 100 57848 400
rect 58464 100 58520 400
rect 59136 100 59192 400
rect 59808 100 59864 400
<< obsm2 >>
rect 14 67930 59850 67970
rect 86 67570 642 67930
rect 758 67570 1314 67930
rect 1430 67570 1986 67930
rect 2102 67570 2658 67930
rect 2774 67570 3330 67930
rect 3446 67570 3666 67930
rect 3782 67570 4338 67930
rect 4454 67570 5010 67930
rect 5126 67570 5682 67930
rect 5798 67570 6354 67930
rect 6470 67570 7026 67930
rect 7142 67570 7362 67930
rect 7478 67570 8034 67930
rect 8150 67570 8706 67930
rect 8822 67570 9378 67930
rect 9494 67570 10050 67930
rect 10166 67570 10722 67930
rect 10838 67570 11058 67930
rect 11174 67570 11730 67930
rect 11846 67570 12402 67930
rect 12518 67570 13074 67930
rect 13190 67570 13746 67930
rect 13862 67570 14418 67930
rect 14534 67570 14754 67930
rect 14870 67570 15426 67930
rect 15542 67570 16098 67930
rect 16214 67570 16770 67930
rect 16886 67570 17442 67930
rect 17558 67570 18114 67930
rect 18230 67570 18450 67930
rect 18566 67570 19122 67930
rect 19238 67570 19794 67930
rect 19910 67570 20466 67930
rect 20582 67570 21138 67930
rect 21254 67570 21810 67930
rect 21926 67570 22146 67930
rect 22262 67570 22818 67930
rect 22934 67570 23490 67930
rect 23606 67570 24162 67930
rect 24278 67570 24834 67930
rect 24950 67570 25506 67930
rect 25622 67570 25842 67930
rect 25958 67570 26514 67930
rect 26630 67570 27186 67930
rect 27302 67570 27858 67930
rect 27974 67570 28530 67930
rect 28646 67570 29202 67930
rect 29318 67570 29874 67930
rect 29990 67570 30210 67930
rect 30326 67570 30882 67930
rect 30998 67570 31554 67930
rect 31670 67570 32226 67930
rect 32342 67570 32898 67930
rect 33014 67570 33570 67930
rect 33686 67570 33906 67930
rect 34022 67570 34578 67930
rect 34694 67570 35250 67930
rect 35366 67570 35922 67930
rect 36038 67570 36594 67930
rect 36710 67570 37266 67930
rect 37382 67570 37602 67930
rect 37718 67570 38274 67930
rect 38390 67570 38946 67930
rect 39062 67570 39618 67930
rect 39734 67570 40290 67930
rect 40406 67570 40962 67930
rect 41078 67570 41298 67930
rect 41414 67570 41970 67930
rect 42086 67570 42642 67930
rect 42758 67570 43314 67930
rect 43430 67570 43986 67930
rect 44102 67570 44658 67930
rect 44774 67570 44994 67930
rect 45110 67570 45666 67930
rect 45782 67570 46338 67930
rect 46454 67570 47010 67930
rect 47126 67570 47682 67930
rect 47798 67570 48354 67930
rect 48470 67570 48690 67930
rect 48806 67570 49362 67930
rect 49478 67570 50034 67930
rect 50150 67570 50706 67930
rect 50822 67570 51378 67930
rect 51494 67570 52050 67930
rect 52166 67570 52386 67930
rect 52502 67570 53058 67930
rect 53174 67570 53730 67930
rect 53846 67570 54402 67930
rect 54518 67570 55074 67930
rect 55190 67570 55746 67930
rect 55862 67570 56082 67930
rect 56198 67570 56754 67930
rect 56870 67570 57426 67930
rect 57542 67570 58098 67930
rect 58214 67570 58770 67930
rect 58886 67570 59442 67930
rect 59558 67570 59778 67930
rect 14 430 59850 67570
rect 86 70 306 430
rect 422 70 978 430
rect 1094 70 1650 430
rect 1766 70 2322 430
rect 2438 70 2994 430
rect 3110 70 3666 430
rect 3782 70 4002 430
rect 4118 70 4674 430
rect 4790 70 5346 430
rect 5462 70 6018 430
rect 6134 70 6690 430
rect 6806 70 7362 430
rect 7478 70 7698 430
rect 7814 70 8370 430
rect 8486 70 9042 430
rect 9158 70 9714 430
rect 9830 70 10386 430
rect 10502 70 11058 430
rect 11174 70 11394 430
rect 11510 70 12066 430
rect 12182 70 12738 430
rect 12854 70 13410 430
rect 13526 70 14082 430
rect 14198 70 14754 430
rect 14870 70 15090 430
rect 15206 70 15762 430
rect 15878 70 16434 430
rect 16550 70 17106 430
rect 17222 70 17778 430
rect 17894 70 18450 430
rect 18566 70 18786 430
rect 18902 70 19458 430
rect 19574 70 20130 430
rect 20246 70 20802 430
rect 20918 70 21474 430
rect 21590 70 22146 430
rect 22262 70 22482 430
rect 22598 70 23154 430
rect 23270 70 23826 430
rect 23942 70 24498 430
rect 24614 70 25170 430
rect 25286 70 25842 430
rect 25958 70 26178 430
rect 26294 70 26850 430
rect 26966 70 27522 430
rect 27638 70 28194 430
rect 28310 70 28866 430
rect 28982 70 29538 430
rect 29654 70 29874 430
rect 29990 70 30546 430
rect 30662 70 31218 430
rect 31334 70 31890 430
rect 32006 70 32562 430
rect 32678 70 33234 430
rect 33350 70 33906 430
rect 34022 70 34242 430
rect 34358 70 34914 430
rect 35030 70 35586 430
rect 35702 70 36258 430
rect 36374 70 36930 430
rect 37046 70 37602 430
rect 37718 70 37938 430
rect 38054 70 38610 430
rect 38726 70 39282 430
rect 39398 70 39954 430
rect 40070 70 40626 430
rect 40742 70 41298 430
rect 41414 70 41634 430
rect 41750 70 42306 430
rect 42422 70 42978 430
rect 43094 70 43650 430
rect 43766 70 44322 430
rect 44438 70 44994 430
rect 45110 70 45330 430
rect 45446 70 46002 430
rect 46118 70 46674 430
rect 46790 70 47346 430
rect 47462 70 48018 430
rect 48134 70 48690 430
rect 48806 70 49026 430
rect 49142 70 49698 430
rect 49814 70 50370 430
rect 50486 70 51042 430
rect 51158 70 51714 430
rect 51830 70 52386 430
rect 52502 70 52722 430
rect 52838 70 53394 430
rect 53510 70 54066 430
rect 54182 70 54738 430
rect 54854 70 55410 430
rect 55526 70 56082 430
rect 56198 70 56418 430
rect 56534 70 57090 430
rect 57206 70 57762 430
rect 57878 70 58434 430
rect 58550 70 59106 430
rect 59222 70 59778 430
rect 14 9 59850 70
<< metal3 >>
rect 100 67872 400 67928
rect 59600 67536 59900 67592
rect 100 67200 400 67256
rect 59600 66864 59900 66920
rect 100 66528 400 66584
rect 59600 66192 59900 66248
rect 100 65856 400 65912
rect 59600 65520 59900 65576
rect 100 65184 400 65240
rect 59600 64848 59900 64904
rect 100 64512 400 64568
rect 59600 64176 59900 64232
rect 100 63840 400 63896
rect 59600 63840 59900 63896
rect 100 63504 400 63560
rect 59600 63168 59900 63224
rect 100 62832 400 62888
rect 59600 62496 59900 62552
rect 100 62160 400 62216
rect 59600 61824 59900 61880
rect 100 61488 400 61544
rect 59600 61152 59900 61208
rect 100 60816 400 60872
rect 59600 60480 59900 60536
rect 100 60144 400 60200
rect 59600 60144 59900 60200
rect 100 59808 400 59864
rect 59600 59472 59900 59528
rect 100 59136 400 59192
rect 59600 58800 59900 58856
rect 100 58464 400 58520
rect 59600 58128 59900 58184
rect 100 57792 400 57848
rect 59600 57456 59900 57512
rect 100 57120 400 57176
rect 59600 56784 59900 56840
rect 100 56448 400 56504
rect 59600 56448 59900 56504
rect 100 56112 400 56168
rect 59600 55776 59900 55832
rect 100 55440 400 55496
rect 59600 55104 59900 55160
rect 100 54768 400 54824
rect 59600 54432 59900 54488
rect 100 54096 400 54152
rect 59600 53760 59900 53816
rect 100 53424 400 53480
rect 59600 53088 59900 53144
rect 100 52752 400 52808
rect 59600 52752 59900 52808
rect 100 52416 400 52472
rect 59600 52080 59900 52136
rect 100 51744 400 51800
rect 59600 51408 59900 51464
rect 100 51072 400 51128
rect 59600 50736 59900 50792
rect 100 50400 400 50456
rect 59600 50064 59900 50120
rect 100 49728 400 49784
rect 59600 49392 59900 49448
rect 100 49056 400 49112
rect 59600 49056 59900 49112
rect 100 48720 400 48776
rect 59600 48384 59900 48440
rect 100 48048 400 48104
rect 59600 47712 59900 47768
rect 100 47376 400 47432
rect 59600 47040 59900 47096
rect 100 46704 400 46760
rect 59600 46368 59900 46424
rect 100 46032 400 46088
rect 59600 45696 59900 45752
rect 100 45360 400 45416
rect 59600 45360 59900 45416
rect 100 45024 400 45080
rect 59600 44688 59900 44744
rect 100 44352 400 44408
rect 59600 44016 59900 44072
rect 100 43680 400 43736
rect 59600 43344 59900 43400
rect 100 43008 400 43064
rect 59600 42672 59900 42728
rect 100 42336 400 42392
rect 59600 42000 59900 42056
rect 100 41664 400 41720
rect 59600 41664 59900 41720
rect 100 41328 400 41384
rect 59600 40992 59900 41048
rect 100 40656 400 40712
rect 59600 40320 59900 40376
rect 100 39984 400 40040
rect 59600 39648 59900 39704
rect 100 39312 400 39368
rect 59600 38976 59900 39032
rect 100 38640 400 38696
rect 59600 38304 59900 38360
rect 100 37968 400 38024
rect 59600 37968 59900 38024
rect 100 37632 400 37688
rect 59600 37296 59900 37352
rect 100 36960 400 37016
rect 59600 36624 59900 36680
rect 100 36288 400 36344
rect 59600 35952 59900 36008
rect 100 35616 400 35672
rect 59600 35280 59900 35336
rect 100 34944 400 35000
rect 59600 34608 59900 34664
rect 100 34272 400 34328
rect 100 33936 400 33992
rect 59600 33936 59900 33992
rect 59600 33600 59900 33656
rect 100 33264 400 33320
rect 59600 32928 59900 32984
rect 100 32592 400 32648
rect 59600 32256 59900 32312
rect 100 31920 400 31976
rect 59600 31584 59900 31640
rect 100 31248 400 31304
rect 59600 30912 59900 30968
rect 100 30576 400 30632
rect 59600 30240 59900 30296
rect 100 29904 400 29960
rect 59600 29904 59900 29960
rect 100 29568 400 29624
rect 59600 29232 59900 29288
rect 100 28896 400 28952
rect 59600 28560 59900 28616
rect 100 28224 400 28280
rect 59600 27888 59900 27944
rect 100 27552 400 27608
rect 59600 27216 59900 27272
rect 100 26880 400 26936
rect 59600 26544 59900 26600
rect 100 26208 400 26264
rect 59600 26208 59900 26264
rect 100 25872 400 25928
rect 59600 25536 59900 25592
rect 100 25200 400 25256
rect 59600 24864 59900 24920
rect 100 24528 400 24584
rect 59600 24192 59900 24248
rect 100 23856 400 23912
rect 59600 23520 59900 23576
rect 100 23184 400 23240
rect 59600 22848 59900 22904
rect 100 22512 400 22568
rect 59600 22512 59900 22568
rect 100 22176 400 22232
rect 59600 21840 59900 21896
rect 100 21504 400 21560
rect 59600 21168 59900 21224
rect 100 20832 400 20888
rect 59600 20496 59900 20552
rect 100 20160 400 20216
rect 59600 19824 59900 19880
rect 100 19488 400 19544
rect 59600 19152 59900 19208
rect 100 18816 400 18872
rect 59600 18816 59900 18872
rect 100 18480 400 18536
rect 59600 18144 59900 18200
rect 100 17808 400 17864
rect 59600 17472 59900 17528
rect 100 17136 400 17192
rect 59600 16800 59900 16856
rect 100 16464 400 16520
rect 59600 16128 59900 16184
rect 100 15792 400 15848
rect 59600 15456 59900 15512
rect 100 15120 400 15176
rect 59600 15120 59900 15176
rect 100 14784 400 14840
rect 59600 14448 59900 14504
rect 100 14112 400 14168
rect 59600 13776 59900 13832
rect 100 13440 400 13496
rect 59600 13104 59900 13160
rect 100 12768 400 12824
rect 59600 12432 59900 12488
rect 100 12096 400 12152
rect 59600 11760 59900 11816
rect 100 11424 400 11480
rect 59600 11424 59900 11480
rect 100 11088 400 11144
rect 59600 10752 59900 10808
rect 100 10416 400 10472
rect 59600 10080 59900 10136
rect 100 9744 400 9800
rect 59600 9408 59900 9464
rect 100 9072 400 9128
rect 59600 8736 59900 8792
rect 100 8400 400 8456
rect 59600 8064 59900 8120
rect 100 7728 400 7784
rect 59600 7728 59900 7784
rect 100 7392 400 7448
rect 59600 7056 59900 7112
rect 100 6720 400 6776
rect 59600 6384 59900 6440
rect 100 6048 400 6104
rect 59600 5712 59900 5768
rect 100 5376 400 5432
rect 59600 5040 59900 5096
rect 100 4704 400 4760
rect 59600 4368 59900 4424
rect 100 4032 400 4088
rect 59600 4032 59900 4088
rect 100 3696 400 3752
rect 59600 3360 59900 3416
rect 100 3024 400 3080
rect 59600 2688 59900 2744
rect 100 2352 400 2408
rect 59600 2016 59900 2072
rect 100 1680 400 1736
rect 59600 1344 59900 1400
rect 100 1008 400 1064
rect 59600 672 59900 728
rect 100 336 400 392
rect 59600 0 59900 56
<< obsm3 >>
rect 9 67170 70 67242
rect 430 67170 59855 67242
rect 9 66950 59855 67170
rect 9 66834 59570 66950
rect 9 66614 59855 66834
rect 9 66498 70 66614
rect 430 66498 59855 66614
rect 9 66278 59855 66498
rect 9 66162 59570 66278
rect 9 65942 59855 66162
rect 9 65826 70 65942
rect 430 65826 59855 65942
rect 9 65606 59855 65826
rect 9 65490 59570 65606
rect 9 65270 59855 65490
rect 9 65154 70 65270
rect 430 65154 59855 65270
rect 9 64934 59855 65154
rect 9 64818 59570 64934
rect 9 64598 59855 64818
rect 9 64482 70 64598
rect 430 64482 59855 64598
rect 9 64262 59855 64482
rect 9 64146 59570 64262
rect 9 63926 59855 64146
rect 9 63810 70 63926
rect 430 63810 59570 63926
rect 9 63590 59855 63810
rect 9 63474 70 63590
rect 430 63474 59855 63590
rect 9 63254 59855 63474
rect 9 63138 59570 63254
rect 9 62918 59855 63138
rect 9 62802 70 62918
rect 430 62802 59855 62918
rect 9 62582 59855 62802
rect 9 62466 59570 62582
rect 9 62246 59855 62466
rect 9 62130 70 62246
rect 430 62130 59855 62246
rect 9 61910 59855 62130
rect 9 61794 59570 61910
rect 9 61574 59855 61794
rect 9 61458 70 61574
rect 430 61458 59855 61574
rect 9 61238 59855 61458
rect 9 61122 59570 61238
rect 9 60902 59855 61122
rect 9 60786 70 60902
rect 430 60786 59855 60902
rect 9 60566 59855 60786
rect 9 60450 59570 60566
rect 9 60230 59855 60450
rect 9 60114 70 60230
rect 430 60114 59570 60230
rect 9 59894 59855 60114
rect 9 59778 70 59894
rect 430 59778 59855 59894
rect 9 59558 59855 59778
rect 9 59442 59570 59558
rect 9 59222 59855 59442
rect 9 59106 70 59222
rect 430 59106 59855 59222
rect 9 58886 59855 59106
rect 9 58770 59570 58886
rect 9 58550 59855 58770
rect 9 58434 70 58550
rect 430 58434 59855 58550
rect 9 58214 59855 58434
rect 9 58098 59570 58214
rect 9 57878 59855 58098
rect 9 57762 70 57878
rect 430 57762 59855 57878
rect 9 57542 59855 57762
rect 9 57426 59570 57542
rect 9 57206 59855 57426
rect 9 57090 70 57206
rect 430 57090 59855 57206
rect 9 56870 59855 57090
rect 9 56754 59570 56870
rect 9 56534 59855 56754
rect 9 56418 70 56534
rect 430 56418 59570 56534
rect 9 56198 59855 56418
rect 9 56082 70 56198
rect 430 56082 59855 56198
rect 9 55862 59855 56082
rect 9 55746 59570 55862
rect 9 55526 59855 55746
rect 9 55410 70 55526
rect 430 55410 59855 55526
rect 9 55190 59855 55410
rect 9 55074 59570 55190
rect 9 54854 59855 55074
rect 9 54738 70 54854
rect 430 54738 59855 54854
rect 9 54518 59855 54738
rect 9 54402 59570 54518
rect 9 54182 59855 54402
rect 9 54066 70 54182
rect 430 54066 59855 54182
rect 9 53846 59855 54066
rect 9 53730 59570 53846
rect 9 53510 59855 53730
rect 9 53394 70 53510
rect 430 53394 59855 53510
rect 9 53174 59855 53394
rect 9 53058 59570 53174
rect 9 52838 59855 53058
rect 9 52722 70 52838
rect 430 52722 59570 52838
rect 9 52502 59855 52722
rect 9 52386 70 52502
rect 430 52386 59855 52502
rect 9 52166 59855 52386
rect 9 52050 59570 52166
rect 9 51830 59855 52050
rect 9 51714 70 51830
rect 430 51714 59855 51830
rect 9 51494 59855 51714
rect 9 51378 59570 51494
rect 9 51158 59855 51378
rect 9 51042 70 51158
rect 430 51042 59855 51158
rect 9 50822 59855 51042
rect 9 50706 59570 50822
rect 9 50486 59855 50706
rect 9 50370 70 50486
rect 430 50370 59855 50486
rect 9 50150 59855 50370
rect 9 50034 59570 50150
rect 9 49814 59855 50034
rect 9 49698 70 49814
rect 430 49698 59855 49814
rect 9 49478 59855 49698
rect 9 49362 59570 49478
rect 9 49142 59855 49362
rect 9 49026 70 49142
rect 430 49026 59570 49142
rect 9 48806 59855 49026
rect 9 48690 70 48806
rect 430 48690 59855 48806
rect 9 48470 59855 48690
rect 9 48354 59570 48470
rect 9 48134 59855 48354
rect 9 48018 70 48134
rect 430 48018 59855 48134
rect 9 47798 59855 48018
rect 9 47682 59570 47798
rect 9 47462 59855 47682
rect 9 47346 70 47462
rect 430 47346 59855 47462
rect 9 47126 59855 47346
rect 9 47010 59570 47126
rect 9 46790 59855 47010
rect 9 46674 70 46790
rect 430 46674 59855 46790
rect 9 46454 59855 46674
rect 9 46338 59570 46454
rect 9 46118 59855 46338
rect 9 46002 70 46118
rect 430 46002 59855 46118
rect 9 45782 59855 46002
rect 9 45666 59570 45782
rect 9 45446 59855 45666
rect 9 45330 70 45446
rect 430 45330 59570 45446
rect 9 45110 59855 45330
rect 9 44994 70 45110
rect 430 44994 59855 45110
rect 9 44774 59855 44994
rect 9 44658 59570 44774
rect 9 44438 59855 44658
rect 9 44322 70 44438
rect 430 44322 59855 44438
rect 9 44102 59855 44322
rect 9 43986 59570 44102
rect 9 43766 59855 43986
rect 9 43650 70 43766
rect 430 43650 59855 43766
rect 9 43430 59855 43650
rect 9 43314 59570 43430
rect 9 43094 59855 43314
rect 9 42978 70 43094
rect 430 42978 59855 43094
rect 9 42758 59855 42978
rect 9 42642 59570 42758
rect 9 42422 59855 42642
rect 9 42306 70 42422
rect 430 42306 59855 42422
rect 9 42086 59855 42306
rect 9 41970 59570 42086
rect 9 41750 59855 41970
rect 9 41634 70 41750
rect 430 41634 59570 41750
rect 9 41414 59855 41634
rect 9 41298 70 41414
rect 430 41298 59855 41414
rect 9 41078 59855 41298
rect 9 40962 59570 41078
rect 9 40742 59855 40962
rect 9 40626 70 40742
rect 430 40626 59855 40742
rect 9 40406 59855 40626
rect 9 40290 59570 40406
rect 9 40070 59855 40290
rect 9 39954 70 40070
rect 430 39954 59855 40070
rect 9 39734 59855 39954
rect 9 39618 59570 39734
rect 9 39398 59855 39618
rect 9 39282 70 39398
rect 430 39282 59855 39398
rect 9 39062 59855 39282
rect 9 38946 59570 39062
rect 9 38726 59855 38946
rect 9 38610 70 38726
rect 430 38610 59855 38726
rect 9 38390 59855 38610
rect 9 38274 59570 38390
rect 9 38054 59855 38274
rect 9 37938 70 38054
rect 430 37938 59570 38054
rect 9 37718 59855 37938
rect 9 37602 70 37718
rect 430 37602 59855 37718
rect 9 37382 59855 37602
rect 9 37266 59570 37382
rect 9 37046 59855 37266
rect 9 36930 70 37046
rect 430 36930 59855 37046
rect 9 36710 59855 36930
rect 9 36594 59570 36710
rect 9 36374 59855 36594
rect 9 36258 70 36374
rect 430 36258 59855 36374
rect 9 36038 59855 36258
rect 9 35922 59570 36038
rect 9 35702 59855 35922
rect 9 35586 70 35702
rect 430 35586 59855 35702
rect 9 35366 59855 35586
rect 9 35250 59570 35366
rect 9 35030 59855 35250
rect 9 34914 70 35030
rect 430 34914 59855 35030
rect 9 34694 59855 34914
rect 9 34578 59570 34694
rect 9 34358 59855 34578
rect 9 34242 70 34358
rect 430 34242 59855 34358
rect 9 34022 59855 34242
rect 9 33906 70 34022
rect 430 33906 59570 34022
rect 9 33686 59855 33906
rect 9 33570 59570 33686
rect 9 33350 59855 33570
rect 9 33234 70 33350
rect 430 33234 59855 33350
rect 9 33014 59855 33234
rect 9 32898 59570 33014
rect 9 32678 59855 32898
rect 9 32562 70 32678
rect 430 32562 59855 32678
rect 9 32342 59855 32562
rect 9 32226 59570 32342
rect 9 32006 59855 32226
rect 9 31890 70 32006
rect 430 31890 59855 32006
rect 9 31670 59855 31890
rect 9 31554 59570 31670
rect 9 31334 59855 31554
rect 9 31218 70 31334
rect 430 31218 59855 31334
rect 9 30998 59855 31218
rect 9 30882 59570 30998
rect 9 30662 59855 30882
rect 9 30546 70 30662
rect 430 30546 59855 30662
rect 9 30326 59855 30546
rect 9 30210 59570 30326
rect 9 29990 59855 30210
rect 9 29874 70 29990
rect 430 29874 59570 29990
rect 9 29654 59855 29874
rect 9 29538 70 29654
rect 430 29538 59855 29654
rect 9 29318 59855 29538
rect 9 29202 59570 29318
rect 9 28982 59855 29202
rect 9 28866 70 28982
rect 430 28866 59855 28982
rect 9 28646 59855 28866
rect 9 28530 59570 28646
rect 9 28310 59855 28530
rect 9 28194 70 28310
rect 430 28194 59855 28310
rect 9 27974 59855 28194
rect 9 27858 59570 27974
rect 9 27638 59855 27858
rect 9 27522 70 27638
rect 430 27522 59855 27638
rect 9 27302 59855 27522
rect 9 27186 59570 27302
rect 9 26966 59855 27186
rect 9 26850 70 26966
rect 430 26850 59855 26966
rect 9 26630 59855 26850
rect 9 26514 59570 26630
rect 9 26294 59855 26514
rect 9 26178 70 26294
rect 430 26178 59570 26294
rect 9 25958 59855 26178
rect 9 25842 70 25958
rect 430 25842 59855 25958
rect 9 25622 59855 25842
rect 9 25506 59570 25622
rect 9 25286 59855 25506
rect 9 25170 70 25286
rect 430 25170 59855 25286
rect 9 24950 59855 25170
rect 9 24834 59570 24950
rect 9 24614 59855 24834
rect 9 24498 70 24614
rect 430 24498 59855 24614
rect 9 24278 59855 24498
rect 9 24162 59570 24278
rect 9 23942 59855 24162
rect 9 23826 70 23942
rect 430 23826 59855 23942
rect 9 23606 59855 23826
rect 9 23490 59570 23606
rect 9 23270 59855 23490
rect 9 23154 70 23270
rect 430 23154 59855 23270
rect 9 22934 59855 23154
rect 9 22818 59570 22934
rect 9 22598 59855 22818
rect 9 22482 70 22598
rect 430 22482 59570 22598
rect 9 22262 59855 22482
rect 9 22146 70 22262
rect 430 22146 59855 22262
rect 9 21926 59855 22146
rect 9 21810 59570 21926
rect 9 21590 59855 21810
rect 9 21474 70 21590
rect 430 21474 59855 21590
rect 9 21254 59855 21474
rect 9 21138 59570 21254
rect 9 20918 59855 21138
rect 9 20802 70 20918
rect 430 20802 59855 20918
rect 9 20582 59855 20802
rect 9 20466 59570 20582
rect 9 20246 59855 20466
rect 9 20130 70 20246
rect 430 20130 59855 20246
rect 9 19910 59855 20130
rect 9 19794 59570 19910
rect 9 19574 59855 19794
rect 9 19458 70 19574
rect 430 19458 59855 19574
rect 9 19238 59855 19458
rect 9 19122 59570 19238
rect 9 18902 59855 19122
rect 9 18786 70 18902
rect 430 18786 59570 18902
rect 9 18566 59855 18786
rect 9 18450 70 18566
rect 430 18450 59855 18566
rect 9 18230 59855 18450
rect 9 18114 59570 18230
rect 9 17894 59855 18114
rect 9 17778 70 17894
rect 430 17778 59855 17894
rect 9 17558 59855 17778
rect 9 17442 59570 17558
rect 9 17222 59855 17442
rect 9 17106 70 17222
rect 430 17106 59855 17222
rect 9 16886 59855 17106
rect 9 16770 59570 16886
rect 9 16550 59855 16770
rect 9 16434 70 16550
rect 430 16434 59855 16550
rect 9 16214 59855 16434
rect 9 16098 59570 16214
rect 9 15878 59855 16098
rect 9 15762 70 15878
rect 430 15762 59855 15878
rect 9 15542 59855 15762
rect 9 15426 59570 15542
rect 9 15206 59855 15426
rect 9 15090 70 15206
rect 430 15090 59570 15206
rect 9 14870 59855 15090
rect 9 14754 70 14870
rect 430 14754 59855 14870
rect 9 14534 59855 14754
rect 9 14418 59570 14534
rect 9 14198 59855 14418
rect 9 14082 70 14198
rect 430 14082 59855 14198
rect 9 13862 59855 14082
rect 9 13746 59570 13862
rect 9 13526 59855 13746
rect 9 13410 70 13526
rect 430 13410 59855 13526
rect 9 13190 59855 13410
rect 9 13074 59570 13190
rect 9 12854 59855 13074
rect 9 12738 70 12854
rect 430 12738 59855 12854
rect 9 12518 59855 12738
rect 9 12402 59570 12518
rect 9 12182 59855 12402
rect 9 12066 70 12182
rect 430 12066 59855 12182
rect 9 11846 59855 12066
rect 9 11730 59570 11846
rect 9 11510 59855 11730
rect 9 11394 70 11510
rect 430 11394 59570 11510
rect 9 11174 59855 11394
rect 9 11058 70 11174
rect 430 11058 59855 11174
rect 9 10838 59855 11058
rect 9 10722 59570 10838
rect 9 10502 59855 10722
rect 9 10386 70 10502
rect 430 10386 59855 10502
rect 9 10166 59855 10386
rect 9 10050 59570 10166
rect 9 9830 59855 10050
rect 9 9714 70 9830
rect 430 9714 59855 9830
rect 9 9494 59855 9714
rect 9 9378 59570 9494
rect 9 9158 59855 9378
rect 9 9042 70 9158
rect 430 9042 59855 9158
rect 9 8822 59855 9042
rect 9 8706 59570 8822
rect 9 8486 59855 8706
rect 9 8370 70 8486
rect 430 8370 59855 8486
rect 9 8150 59855 8370
rect 9 8034 59570 8150
rect 9 7814 59855 8034
rect 9 7698 70 7814
rect 430 7698 59570 7814
rect 9 7478 59855 7698
rect 9 7362 70 7478
rect 430 7362 59855 7478
rect 9 7142 59855 7362
rect 9 7026 59570 7142
rect 9 6806 59855 7026
rect 9 6690 70 6806
rect 430 6690 59855 6806
rect 9 6470 59855 6690
rect 9 6354 59570 6470
rect 9 6134 59855 6354
rect 9 6018 70 6134
rect 430 6018 59855 6134
rect 9 5798 59855 6018
rect 9 5682 59570 5798
rect 9 5462 59855 5682
rect 9 5346 70 5462
rect 430 5346 59855 5462
rect 9 5126 59855 5346
rect 9 5010 59570 5126
rect 9 4790 59855 5010
rect 9 4674 70 4790
rect 430 4674 59855 4790
rect 9 4454 59855 4674
rect 9 4338 59570 4454
rect 9 4118 59855 4338
rect 9 4002 70 4118
rect 430 4002 59570 4118
rect 9 3782 59855 4002
rect 9 3666 70 3782
rect 430 3666 59855 3782
rect 9 3446 59855 3666
rect 9 3330 59570 3446
rect 9 3110 59855 3330
rect 9 2994 70 3110
rect 430 2994 59855 3110
rect 9 2774 59855 2994
rect 9 2658 59570 2774
rect 9 2438 59855 2658
rect 9 2322 70 2438
rect 430 2322 59855 2438
rect 9 2102 59855 2322
rect 9 1986 59570 2102
rect 9 1766 59855 1986
rect 9 1650 70 1766
rect 430 1650 59855 1766
rect 9 1430 59855 1650
rect 9 1314 59570 1430
rect 9 1094 59855 1314
rect 9 978 70 1094
rect 430 978 59855 1094
rect 9 758 59855 978
rect 9 642 59570 758
rect 9 422 59855 642
rect 9 306 70 422
rect 430 306 59855 422
rect 9 86 59855 306
rect 9 14 59570 86
<< metal4 >>
rect 2224 1538 2384 66278
rect 9904 1538 10064 66278
rect 17584 1538 17744 66278
rect 25264 1538 25424 66278
rect 32944 1538 33104 66278
rect 40624 1538 40784 66278
rect 48304 1538 48464 66278
rect 55984 1538 56144 66278
<< labels >>
rlabel metal3 s 100 44352 400 44408 6 io_in[0]
port 1 nsew signal input
rlabel metal3 s 100 45024 400 45080 6 io_in[10]
port 2 nsew signal input
rlabel metal3 s 100 22176 400 22232 6 io_in[11]
port 3 nsew signal input
rlabel metal3 s 100 38640 400 38696 6 io_in[12]
port 4 nsew signal input
rlabel metal3 s 100 26208 400 26264 6 io_in[13]
port 5 nsew signal input
rlabel metal3 s 100 22512 400 22568 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 29904 67600 29960 67900 6 io_in[15]
port 7 nsew signal input
rlabel metal3 s 59600 16800 59900 16856 6 io_in[16]
port 8 nsew signal input
rlabel metal3 s 59600 64176 59900 64232 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 38976 67600 39032 67900 6 io_in[18]
port 10 nsew signal input
rlabel metal3 s 59600 2688 59900 2744 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 3696 67600 3752 67900 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 47040 67600 47096 67900 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 45024 100 45080 400 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 59808 67600 59864 67900 6 io_in[22]
port 15 nsew signal input
rlabel metal3 s 59600 59472 59900 59528 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 52752 100 52808 400 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 8400 100 8456 400 6 io_in[25]
port 18 nsew signal input
rlabel metal3 s 100 53424 400 53480 6 io_in[26]
port 19 nsew signal input
rlabel metal3 s 100 43680 400 43736 6 io_in[27]
port 20 nsew signal input
rlabel metal3 s 100 49728 400 49784 6 io_in[28]
port 21 nsew signal input
rlabel metal3 s 100 39984 400 40040 6 io_in[29]
port 22 nsew signal input
rlabel metal3 s 59600 67536 59900 67592 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 41664 100 41720 400 6 io_in[30]
port 24 nsew signal input
rlabel metal3 s 100 26880 400 26936 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 54096 100 54152 400 6 io_in[32]
port 26 nsew signal input
rlabel metal3 s 100 6720 400 6776 6 io_in[33]
port 27 nsew signal input
rlabel metal3 s 100 57120 400 57176 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 53088 67600 53144 67900 6 io_in[35]
port 29 nsew signal input
rlabel metal3 s 59600 60480 59900 60536 6 io_in[36]
port 30 nsew signal input
rlabel metal3 s 59600 52752 59900 52808 6 io_in[37]
port 31 nsew signal input
rlabel metal3 s 59600 66864 59900 66920 6 io_in[3]
port 32 nsew signal input
rlabel metal3 s 59600 32928 59900 32984 6 io_in[4]
port 33 nsew signal input
rlabel metal3 s 100 12096 400 12152 6 io_in[5]
port 34 nsew signal input
rlabel metal3 s 59600 16128 59900 16184 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 48384 67600 48440 67900 6 io_in[7]
port 36 nsew signal input
rlabel metal3 s 100 29568 400 29624 6 io_in[8]
port 37 nsew signal input
rlabel metal3 s 100 33264 400 33320 6 io_in[9]
port 38 nsew signal input
rlabel metal3 s 59600 49056 59900 49112 6 io_oeb[0]
port 39 nsew signal output
rlabel metal3 s 59600 45360 59900 45416 6 io_oeb[10]
port 40 nsew signal output
rlabel metal3 s 100 66528 400 66584 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 39312 100 39368 400 6 io_oeb[12]
port 42 nsew signal output
rlabel metal3 s 100 16464 400 16520 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 58464 100 58520 400 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 36624 67600 36680 67900 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 18480 100 18536 400 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 6048 100 6104 400 6 io_oeb[17]
port 47 nsew signal output
rlabel metal3 s 100 67200 400 67256 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 18480 67600 18536 67900 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 13104 67600 13160 67900 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 32928 67600 32984 67900 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 54768 100 54824 400 6 io_oeb[21]
port 52 nsew signal output
rlabel metal3 s 59600 20496 59900 20552 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 58128 67600 58184 67900 6 io_oeb[23]
port 54 nsew signal output
rlabel metal3 s 100 18480 400 18536 6 io_oeb[24]
port 55 nsew signal output
rlabel metal3 s 100 9072 400 9128 6 io_oeb[25]
port 56 nsew signal output
rlabel metal3 s 100 58464 400 58520 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 53424 100 53480 400 6 io_oeb[27]
port 58 nsew signal output
rlabel metal3 s 100 65184 400 65240 6 io_oeb[28]
port 59 nsew signal output
rlabel metal3 s 59600 36624 59900 36680 6 io_oeb[29]
port 60 nsew signal output
rlabel metal3 s 59600 28560 59900 28616 6 io_oeb[2]
port 61 nsew signal output
rlabel metal3 s 59600 0 59900 56 6 io_oeb[30]
port 62 nsew signal output
rlabel metal3 s 100 19488 400 19544 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 52080 67600 52136 67900 6 io_oeb[32]
port 64 nsew signal output
rlabel metal3 s 59600 14448 59900 14504 6 io_oeb[33]
port 65 nsew signal output
rlabel metal3 s 100 52416 400 52472 6 io_oeb[34]
port 66 nsew signal output
rlabel metal3 s 59600 61824 59900 61880 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 31584 67600 31640 67900 6 io_oeb[36]
port 68 nsew signal output
rlabel metal3 s 59600 29904 59900 29960 6 io_oeb[37]
port 69 nsew signal output
rlabel metal3 s 100 48048 400 48104 6 io_oeb[3]
port 70 nsew signal output
rlabel metal3 s 100 8400 400 8456 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 42672 67600 42728 67900 6 io_oeb[5]
port 72 nsew signal output
rlabel metal3 s 100 50400 400 50456 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 26544 67600 26600 67900 6 io_oeb[7]
port 74 nsew signal output
rlabel metal3 s 100 31920 400 31976 6 io_oeb[8]
port 75 nsew signal output
rlabel metal3 s 59600 66192 59900 66248 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 6384 67600 6440 67900 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 15456 67600 15512 67900 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 41328 100 41384 400 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 58800 67600 58856 67900 6 io_out[12]
port 80 nsew signal output
rlabel metal3 s 100 63840 400 63896 6 io_out[13]
port 81 nsew signal output
rlabel metal3 s 100 47376 400 47432 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 25872 100 25928 400 6 io_out[15]
port 83 nsew signal output
rlabel metal3 s 59600 57456 59900 57512 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 7392 100 7448 400 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 59808 100 59864 400 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 10080 67600 10136 67900 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 4032 100 4088 400 6 io_out[1]
port 88 nsew signal output
rlabel metal3 s 59600 10080 59900 10136 6 io_out[20]
port 89 nsew signal output
rlabel metal3 s 100 42336 400 42392 6 io_out[21]
port 90 nsew signal output
rlabel metal3 s 59600 18144 59900 18200 6 io_out[22]
port 91 nsew signal output
rlabel metal3 s 100 23856 400 23912 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 56112 100 56168 400 6 io_out[24]
port 93 nsew signal output
rlabel metal3 s 59600 5712 59900 5768 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 26880 100 26936 400 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 21504 100 21560 400 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 40992 67600 41048 67900 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 43680 100 43736 400 6 io_out[29]
port 98 nsew signal output
rlabel metal3 s 59600 26544 59900 26600 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 54432 67600 54488 67900 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 22512 100 22568 400 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 35952 67600 36008 67900 6 io_out[32]
port 102 nsew signal output
rlabel metal3 s 100 23184 400 23240 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 42336 100 42392 400 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 37968 100 38024 400 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 15120 100 15176 400 6 io_out[36]
port 106 nsew signal output
rlabel metal3 s 100 3024 400 3080 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 25536 67600 25592 67900 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 29568 100 29624 400 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 22848 67600 22904 67900 6 io_out[5]
port 110 nsew signal output
rlabel metal3 s 100 11424 400 11480 6 io_out[6]
port 111 nsew signal output
rlabel metal3 s 100 36288 400 36344 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 46704 100 46760 400 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 16464 100 16520 400 6 io_out[9]
port 114 nsew signal output
rlabel metal3 s 100 32592 400 32648 6 la_data_in[0]
port 115 nsew signal input
rlabel metal3 s 59600 63840 59900 63896 6 la_data_in[10]
port 116 nsew signal input
rlabel metal3 s 59600 32256 59900 32312 6 la_data_in[11]
port 117 nsew signal input
rlabel metal2 s 19488 100 19544 400 6 la_data_in[12]
port 118 nsew signal input
rlabel metal2 s 21840 67600 21896 67900 6 la_data_in[13]
port 119 nsew signal input
rlabel metal3 s 100 56112 400 56168 6 la_data_in[14]
port 120 nsew signal input
rlabel metal3 s 59600 50064 59900 50120 6 la_data_in[15]
port 121 nsew signal input
rlabel metal2 s 2016 67600 2072 67900 6 la_data_in[16]
port 122 nsew signal input
rlabel metal3 s 59600 13776 59900 13832 6 la_data_in[17]
port 123 nsew signal input
rlabel metal2 s 27888 67600 27944 67900 6 la_data_in[18]
port 124 nsew signal input
rlabel metal3 s 100 9744 400 9800 6 la_data_in[19]
port 125 nsew signal input
rlabel metal2 s 10752 67600 10808 67900 6 la_data_in[1]
port 126 nsew signal input
rlabel metal3 s 59600 17472 59900 17528 6 la_data_in[20]
port 127 nsew signal input
rlabel metal3 s 100 48720 400 48776 6 la_data_in[21]
port 128 nsew signal input
rlabel metal3 s 100 28224 400 28280 6 la_data_in[22]
port 129 nsew signal input
rlabel metal3 s 59600 52080 59900 52136 6 la_data_in[23]
port 130 nsew signal input
rlabel metal2 s 28560 67600 28616 67900 6 la_data_in[24]
port 131 nsew signal input
rlabel metal2 s 9408 67600 9464 67900 6 la_data_in[25]
port 132 nsew signal input
rlabel metal2 s 35280 67600 35336 67900 6 la_data_in[26]
port 133 nsew signal input
rlabel metal3 s 100 57792 400 57848 6 la_data_in[27]
port 134 nsew signal input
rlabel metal3 s 100 60144 400 60200 6 la_data_in[28]
port 135 nsew signal input
rlabel metal3 s 59600 19824 59900 19880 6 la_data_in[29]
port 136 nsew signal input
rlabel metal2 s 24192 67600 24248 67900 6 la_data_in[2]
port 137 nsew signal input
rlabel metal3 s 100 4704 400 4760 6 la_data_in[30]
port 138 nsew signal input
rlabel metal2 s 50064 67600 50120 67900 6 la_data_in[31]
port 139 nsew signal input
rlabel metal3 s 100 25872 400 25928 6 la_data_in[32]
port 140 nsew signal input
rlabel metal3 s 100 43008 400 43064 6 la_data_in[33]
port 141 nsew signal input
rlabel metal2 s 672 67600 728 67900 6 la_data_in[34]
port 142 nsew signal input
rlabel metal3 s 100 56448 400 56504 6 la_data_in[35]
port 143 nsew signal input
rlabel metal2 s 45360 100 45416 400 6 la_data_in[36]
port 144 nsew signal input
rlabel metal3 s 100 62832 400 62888 6 la_data_in[37]
port 145 nsew signal input
rlabel metal2 s 28896 100 28952 400 6 la_data_in[38]
port 146 nsew signal input
rlabel metal2 s 30912 67600 30968 67900 6 la_data_in[39]
port 147 nsew signal input
rlabel metal3 s 59600 38976 59900 39032 6 la_data_in[3]
port 148 nsew signal input
rlabel metal2 s 22176 100 22232 400 6 la_data_in[40]
port 149 nsew signal input
rlabel metal2 s 30576 100 30632 400 6 la_data_in[41]
port 150 nsew signal input
rlabel metal3 s 100 21504 400 21560 6 la_data_in[42]
port 151 nsew signal input
rlabel metal2 s 56112 67600 56168 67900 6 la_data_in[43]
port 152 nsew signal input
rlabel metal3 s 59600 4368 59900 4424 6 la_data_in[44]
port 153 nsew signal input
rlabel metal2 s 20832 100 20888 400 6 la_data_in[45]
port 154 nsew signal input
rlabel metal3 s 59600 50736 59900 50792 6 la_data_in[46]
port 155 nsew signal input
rlabel metal2 s 39984 100 40040 400 6 la_data_in[47]
port 156 nsew signal input
rlabel metal2 s 25872 67600 25928 67900 6 la_data_in[48]
port 157 nsew signal input
rlabel metal2 s 20496 67600 20552 67900 6 la_data_in[49]
port 158 nsew signal input
rlabel metal2 s 1344 67600 1400 67900 6 la_data_in[4]
port 159 nsew signal input
rlabel metal2 s 21168 67600 21224 67900 6 la_data_in[50]
port 160 nsew signal input
rlabel metal2 s 29904 100 29960 400 6 la_data_in[51]
port 161 nsew signal input
rlabel metal3 s 59600 25536 59900 25592 6 la_data_in[52]
port 162 nsew signal input
rlabel metal2 s 45696 67600 45752 67900 6 la_data_in[53]
port 163 nsew signal input
rlabel metal2 s 41328 67600 41384 67900 6 la_data_in[54]
port 164 nsew signal input
rlabel metal3 s 100 17136 400 17192 6 la_data_in[55]
port 165 nsew signal input
rlabel metal3 s 100 18816 400 18872 6 la_data_in[56]
port 166 nsew signal input
rlabel metal3 s 100 65856 400 65912 6 la_data_in[57]
port 167 nsew signal input
rlabel metal2 s 23184 100 23240 400 6 la_data_in[58]
port 168 nsew signal input
rlabel metal3 s 59600 62496 59900 62552 6 la_data_in[59]
port 169 nsew signal input
rlabel metal2 s 11088 100 11144 400 6 la_data_in[5]
port 170 nsew signal input
rlabel metal3 s 59600 46368 59900 46424 6 la_data_in[60]
port 171 nsew signal input
rlabel metal3 s 100 1680 400 1736 6 la_data_in[61]
port 172 nsew signal input
rlabel metal2 s 37632 100 37688 400 6 la_data_in[62]
port 173 nsew signal input
rlabel metal2 s 12432 67600 12488 67900 6 la_data_in[63]
port 174 nsew signal input
rlabel metal2 s 12768 100 12824 400 6 la_data_in[6]
port 175 nsew signal input
rlabel metal3 s 59600 27216 59900 27272 6 la_data_in[7]
port 176 nsew signal input
rlabel metal3 s 100 1008 400 1064 6 la_data_in[8]
port 177 nsew signal input
rlabel metal2 s 53760 67600 53816 67900 6 la_data_in[9]
port 178 nsew signal input
rlabel metal2 s 51408 67600 51464 67900 6 la_data_out[0]
port 179 nsew signal output
rlabel metal3 s 59600 38304 59900 38360 6 la_data_out[10]
port 180 nsew signal output
rlabel metal3 s 100 2352 400 2408 6 la_data_out[11]
port 181 nsew signal output
rlabel metal3 s 100 46032 400 46088 6 la_data_out[12]
port 182 nsew signal output
rlabel metal2 s 23856 100 23912 400 6 la_data_out[13]
port 183 nsew signal output
rlabel metal3 s 59600 30240 59900 30296 6 la_data_out[14]
port 184 nsew signal output
rlabel metal3 s 100 54768 400 54824 6 la_data_out[15]
port 185 nsew signal output
rlabel metal3 s 59600 39648 59900 39704 6 la_data_out[16]
port 186 nsew signal output
rlabel metal2 s 27216 67600 27272 67900 6 la_data_out[17]
port 187 nsew signal output
rlabel metal3 s 59600 56784 59900 56840 6 la_data_out[18]
port 188 nsew signal output
rlabel metal2 s 33936 100 33992 400 6 la_data_out[19]
port 189 nsew signal output
rlabel metal3 s 59600 33936 59900 33992 6 la_data_out[1]
port 190 nsew signal output
rlabel metal3 s 59600 13104 59900 13160 6 la_data_out[20]
port 191 nsew signal output
rlabel metal3 s 100 63504 400 63560 6 la_data_out[21]
port 192 nsew signal output
rlabel metal3 s 59600 44016 59900 44072 6 la_data_out[22]
port 193 nsew signal output
rlabel metal2 s 18816 100 18872 400 6 la_data_out[23]
port 194 nsew signal output
rlabel metal3 s 100 28896 400 28952 6 la_data_out[24]
port 195 nsew signal output
rlabel metal2 s 34272 100 34328 400 6 la_data_out[25]
port 196 nsew signal output
rlabel metal3 s 100 62160 400 62216 6 la_data_out[26]
port 197 nsew signal output
rlabel metal2 s 34608 67600 34664 67900 6 la_data_out[27]
port 198 nsew signal output
rlabel metal3 s 59600 55104 59900 55160 6 la_data_out[28]
port 199 nsew signal output
rlabel metal2 s 27552 100 27608 400 6 la_data_out[29]
port 200 nsew signal output
rlabel metal3 s 100 14784 400 14840 6 la_data_out[2]
port 201 nsew signal output
rlabel metal3 s 59600 33600 59900 33656 6 la_data_out[30]
port 202 nsew signal output
rlabel metal3 s 59600 7056 59900 7112 6 la_data_out[31]
port 203 nsew signal output
rlabel metal2 s 33600 67600 33656 67900 6 la_data_out[32]
port 204 nsew signal output
rlabel metal3 s 59600 15456 59900 15512 6 la_data_out[33]
port 205 nsew signal output
rlabel metal2 s 31248 100 31304 400 6 la_data_out[34]
port 206 nsew signal output
rlabel metal2 s 30240 67600 30296 67900 6 la_data_out[35]
port 207 nsew signal output
rlabel metal3 s 59600 55776 59900 55832 6 la_data_out[36]
port 208 nsew signal output
rlabel metal3 s 59600 29232 59900 29288 6 la_data_out[37]
port 209 nsew signal output
rlabel metal3 s 59600 5040 59900 5096 6 la_data_out[38]
port 210 nsew signal output
rlabel metal3 s 59600 12432 59900 12488 6 la_data_out[39]
port 211 nsew signal output
rlabel metal3 s 100 10416 400 10472 6 la_data_out[3]
port 212 nsew signal output
rlabel metal3 s 59600 2016 59900 2072 6 la_data_out[40]
port 213 nsew signal output
rlabel metal3 s 59600 23520 59900 23576 6 la_data_out[41]
port 214 nsew signal output
rlabel metal3 s 59600 58128 59900 58184 6 la_data_out[42]
port 215 nsew signal output
rlabel metal2 s 3696 100 3752 400 6 la_data_out[43]
port 216 nsew signal output
rlabel metal2 s 26208 100 26264 400 6 la_data_out[44]
port 217 nsew signal output
rlabel metal2 s 5712 67600 5768 67900 6 la_data_out[45]
port 218 nsew signal output
rlabel metal2 s 5040 67600 5096 67900 6 la_data_out[46]
port 219 nsew signal output
rlabel metal3 s 100 45360 400 45416 6 la_data_out[47]
port 220 nsew signal output
rlabel metal2 s 14784 100 14840 400 6 la_data_out[48]
port 221 nsew signal output
rlabel metal2 s 57792 100 57848 400 6 la_data_out[49]
port 222 nsew signal output
rlabel metal2 s 32256 67600 32312 67900 6 la_data_out[4]
port 223 nsew signal output
rlabel metal2 s 18144 67600 18200 67900 6 la_data_out[50]
port 224 nsew signal output
rlabel metal3 s 100 61488 400 61544 6 la_data_out[51]
port 225 nsew signal output
rlabel metal3 s 59600 8064 59900 8120 6 la_data_out[52]
port 226 nsew signal output
rlabel metal3 s 100 60816 400 60872 6 la_data_out[53]
port 227 nsew signal output
rlabel metal3 s 59600 47712 59900 47768 6 la_data_out[54]
port 228 nsew signal output
rlabel metal2 s 19824 67600 19880 67900 6 la_data_out[55]
port 229 nsew signal output
rlabel metal3 s 59600 19152 59900 19208 6 la_data_out[56]
port 230 nsew signal output
rlabel metal2 s 44688 67600 44744 67900 6 la_data_out[57]
port 231 nsew signal output
rlabel metal3 s 59600 48384 59900 48440 6 la_data_out[58]
port 232 nsew signal output
rlabel metal3 s 100 24528 400 24584 6 la_data_out[59]
port 233 nsew signal output
rlabel metal3 s 59600 42000 59900 42056 6 la_data_out[5]
port 234 nsew signal output
rlabel metal2 s 47712 67600 47768 67900 6 la_data_out[60]
port 235 nsew signal output
rlabel metal2 s 17136 100 17192 400 6 la_data_out[61]
port 236 nsew signal output
rlabel metal2 s 55440 100 55496 400 6 la_data_out[62]
port 237 nsew signal output
rlabel metal3 s 59600 8736 59900 8792 6 la_data_out[63]
port 238 nsew signal output
rlabel metal3 s 59600 22512 59900 22568 6 la_data_out[6]
port 239 nsew signal output
rlabel metal2 s 57456 67600 57512 67900 6 la_data_out[7]
port 240 nsew signal output
rlabel metal3 s 100 3696 400 3752 6 la_data_out[8]
port 241 nsew signal output
rlabel metal3 s 59600 34608 59900 34664 6 la_data_out[9]
port 242 nsew signal output
rlabel metal3 s 59600 27888 59900 27944 6 la_oenb[0]
port 243 nsew signal input
rlabel metal3 s 59600 49392 59900 49448 6 la_oenb[10]
port 244 nsew signal input
rlabel metal3 s 59600 40320 59900 40376 6 la_oenb[11]
port 245 nsew signal input
rlabel metal3 s 100 64512 400 64568 6 la_oenb[12]
port 246 nsew signal input
rlabel metal3 s 100 51072 400 51128 6 la_oenb[13]
port 247 nsew signal input
rlabel metal2 s 47376 100 47432 400 6 la_oenb[14]
port 248 nsew signal input
rlabel metal2 s 56448 100 56504 400 6 la_oenb[15]
port 249 nsew signal input
rlabel metal2 s 9072 100 9128 400 6 la_oenb[16]
port 250 nsew signal input
rlabel metal3 s 100 7728 400 7784 6 la_oenb[17]
port 251 nsew signal input
rlabel metal2 s 0 67600 56 67900 6 la_oenb[18]
port 252 nsew signal input
rlabel metal3 s 59600 9408 59900 9464 6 la_oenb[19]
port 253 nsew signal input
rlabel metal2 s 8064 67600 8120 67900 6 la_oenb[1]
port 254 nsew signal input
rlabel metal3 s 100 37632 400 37688 6 la_oenb[20]
port 255 nsew signal input
rlabel metal2 s 22176 67600 22232 67900 6 la_oenb[21]
port 256 nsew signal input
rlabel metal2 s 43344 67600 43400 67900 6 la_oenb[22]
port 257 nsew signal input
rlabel metal2 s 17808 100 17864 400 6 la_oenb[23]
port 258 nsew signal input
rlabel metal3 s 59600 43344 59900 43400 6 la_oenb[24]
port 259 nsew signal input
rlabel metal2 s 57120 100 57176 400 6 la_oenb[25]
port 260 nsew signal input
rlabel metal2 s 8736 67600 8792 67900 6 la_oenb[26]
port 261 nsew signal input
rlabel metal2 s 11424 100 11480 400 6 la_oenb[27]
port 262 nsew signal input
rlabel metal3 s 100 39312 400 39368 6 la_oenb[28]
port 263 nsew signal input
rlabel metal3 s 59600 64848 59900 64904 6 la_oenb[29]
port 264 nsew signal input
rlabel metal2 s 59472 67600 59528 67900 6 la_oenb[2]
port 265 nsew signal input
rlabel metal3 s 59600 58800 59900 58856 6 la_oenb[30]
port 266 nsew signal input
rlabel metal2 s 23520 67600 23576 67900 6 la_oenb[31]
port 267 nsew signal input
rlabel metal3 s 59600 56448 59900 56504 6 la_oenb[32]
port 268 nsew signal input
rlabel metal2 s 32592 100 32648 400 6 la_oenb[33]
port 269 nsew signal input
rlabel metal2 s 7056 67600 7112 67900 6 la_oenb[34]
port 270 nsew signal input
rlabel metal2 s 1680 100 1736 400 6 la_oenb[35]
port 271 nsew signal input
rlabel metal2 s 336 100 392 400 6 la_oenb[36]
port 272 nsew signal input
rlabel metal2 s 4368 67600 4424 67900 6 la_oenb[37]
port 273 nsew signal input
rlabel metal2 s 33264 100 33320 400 6 la_oenb[38]
port 274 nsew signal input
rlabel metal3 s 100 27552 400 27608 6 la_oenb[39]
port 275 nsew signal input
rlabel metal3 s 100 34944 400 35000 6 la_oenb[3]
port 276 nsew signal input
rlabel metal3 s 59600 11760 59900 11816 6 la_oenb[40]
port 277 nsew signal input
rlabel metal2 s 19152 67600 19208 67900 6 la_oenb[41]
port 278 nsew signal input
rlabel metal3 s 100 40656 400 40712 6 la_oenb[42]
port 279 nsew signal input
rlabel metal2 s 12096 100 12152 400 6 la_oenb[43]
port 280 nsew signal input
rlabel metal2 s 28224 100 28280 400 6 la_oenb[44]
port 281 nsew signal input
rlabel metal2 s 48720 67600 48776 67900 6 la_oenb[45]
port 282 nsew signal input
rlabel metal2 s 51072 100 51128 400 6 la_oenb[46]
port 283 nsew signal input
rlabel metal3 s 100 7392 400 7448 6 la_oenb[47]
port 284 nsew signal input
rlabel metal3 s 100 46704 400 46760 6 la_oenb[48]
port 285 nsew signal input
rlabel metal3 s 100 336 400 392 6 la_oenb[49]
port 286 nsew signal input
rlabel metal3 s 100 59808 400 59864 6 la_oenb[4]
port 287 nsew signal input
rlabel metal2 s 49056 100 49112 400 6 la_oenb[50]
port 288 nsew signal input
rlabel metal2 s 16800 67600 16856 67900 6 la_oenb[51]
port 289 nsew signal input
rlabel metal3 s 59600 3360 59900 3416 6 la_oenb[52]
port 290 nsew signal input
rlabel metal3 s 59600 44688 59900 44744 6 la_oenb[53]
port 291 nsew signal input
rlabel metal3 s 100 34272 400 34328 6 la_oenb[54]
port 292 nsew signal input
rlabel metal3 s 59600 37296 59900 37352 6 la_oenb[55]
port 293 nsew signal input
rlabel metal2 s 48720 100 48776 400 6 la_oenb[56]
port 294 nsew signal input
rlabel metal2 s 52416 67600 52472 67900 6 la_oenb[57]
port 295 nsew signal input
rlabel metal3 s 59600 10752 59900 10808 6 la_oenb[58]
port 296 nsew signal input
rlabel metal2 s 33936 67600 33992 67900 6 la_oenb[59]
port 297 nsew signal input
rlabel metal2 s 59136 100 59192 400 6 la_oenb[5]
port 298 nsew signal input
rlabel metal3 s 100 31248 400 31304 6 la_oenb[60]
port 299 nsew signal input
rlabel metal2 s 7728 100 7784 400 6 la_oenb[61]
port 300 nsew signal input
rlabel metal3 s 59600 35952 59900 36008 6 la_oenb[62]
port 301 nsew signal input
rlabel metal3 s 100 15120 400 15176 6 la_oenb[63]
port 302 nsew signal input
rlabel metal3 s 59600 45696 59900 45752 6 la_oenb[6]
port 303 nsew signal input
rlabel metal2 s 15792 100 15848 400 6 la_oenb[7]
port 304 nsew signal input
rlabel metal3 s 59600 672 59900 728 6 la_oenb[8]
port 305 nsew signal input
rlabel metal2 s 14448 67600 14504 67900 6 la_oenb[9]
port 306 nsew signal input
rlabel metal2 s 50736 67600 50792 67900 6 user_clock2
port 307 nsew signal input
rlabel metal3 s 59600 53088 59900 53144 6 user_irq[0]
port 308 nsew signal output
rlabel metal2 s 11760 67600 11816 67900 6 user_irq[1]
port 309 nsew signal output
rlabel metal3 s 100 41328 400 41384 6 user_irq[2]
port 310 nsew signal output
rlabel metal4 s 2224 1538 2384 66278 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 66278 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 66278 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 48304 1538 48464 66278 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 66278 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 66278 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 40624 1538 40784 66278 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 55984 1538 56144 66278 6 vss
port 312 nsew ground bidirectional
rlabel metal3 s 59600 15120 59900 15176 6 wb_clk_i
port 313 nsew signal input
rlabel metal2 s 7392 67600 7448 67900 6 wb_rst_i
port 314 nsew signal input
rlabel metal3 s 59600 26208 59900 26264 6 wbs_ack_o
port 315 nsew signal output
rlabel metal2 s 38304 67600 38360 67900 6 wbs_adr_i[0]
port 316 nsew signal input
rlabel metal2 s 24864 67600 24920 67900 6 wbs_adr_i[10]
port 317 nsew signal input
rlabel metal3 s 100 36960 400 37016 6 wbs_adr_i[11]
port 318 nsew signal input
rlabel metal2 s 5376 100 5432 400 6 wbs_adr_i[12]
port 319 nsew signal input
rlabel metal2 s 35616 100 35672 400 6 wbs_adr_i[13]
port 320 nsew signal input
rlabel metal3 s 100 6048 400 6104 6 wbs_adr_i[14]
port 321 nsew signal input
rlabel metal3 s 59600 47040 59900 47096 6 wbs_adr_i[15]
port 322 nsew signal input
rlabel metal2 s 40656 100 40712 400 6 wbs_adr_i[16]
port 323 nsew signal input
rlabel metal3 s 100 35616 400 35672 6 wbs_adr_i[17]
port 324 nsew signal input
rlabel metal3 s 59600 24192 59900 24248 6 wbs_adr_i[18]
port 325 nsew signal input
rlabel metal3 s 59600 1344 59900 1400 6 wbs_adr_i[19]
port 326 nsew signal input
rlabel metal3 s 100 4032 400 4088 6 wbs_adr_i[1]
port 327 nsew signal input
rlabel metal2 s 55776 67600 55832 67900 6 wbs_adr_i[20]
port 328 nsew signal input
rlabel metal2 s 36288 100 36344 400 6 wbs_adr_i[21]
port 329 nsew signal input
rlabel metal2 s 51744 100 51800 400 6 wbs_adr_i[22]
port 330 nsew signal input
rlabel metal3 s 59600 18816 59900 18872 6 wbs_adr_i[23]
port 331 nsew signal input
rlabel metal2 s 3360 67600 3416 67900 6 wbs_adr_i[24]
port 332 nsew signal input
rlabel metal3 s 100 11088 400 11144 6 wbs_adr_i[25]
port 333 nsew signal input
rlabel metal2 s 6720 100 6776 400 6 wbs_adr_i[26]
port 334 nsew signal input
rlabel metal2 s 17472 67600 17528 67900 6 wbs_adr_i[27]
port 335 nsew signal input
rlabel metal3 s 59600 41664 59900 41720 6 wbs_adr_i[28]
port 336 nsew signal input
rlabel metal3 s 59600 65520 59900 65576 6 wbs_adr_i[29]
port 337 nsew signal input
rlabel metal2 s 25200 100 25256 400 6 wbs_adr_i[2]
port 338 nsew signal input
rlabel metal3 s 100 25200 400 25256 6 wbs_adr_i[30]
port 339 nsew signal input
rlabel metal3 s 59600 30912 59900 30968 6 wbs_adr_i[31]
port 340 nsew signal input
rlabel metal2 s 49728 100 49784 400 6 wbs_adr_i[3]
port 341 nsew signal input
rlabel metal2 s 45024 67600 45080 67900 6 wbs_adr_i[4]
port 342 nsew signal input
rlabel metal2 s 48048 100 48104 400 6 wbs_adr_i[5]
port 343 nsew signal input
rlabel metal3 s 100 15792 400 15848 6 wbs_adr_i[6]
port 344 nsew signal input
rlabel metal2 s 3024 100 3080 400 6 wbs_adr_i[7]
port 345 nsew signal input
rlabel metal3 s 59600 4032 59900 4088 6 wbs_adr_i[8]
port 346 nsew signal input
rlabel metal3 s 59600 21168 59900 21224 6 wbs_adr_i[9]
port 347 nsew signal input
rlabel metal2 s 16128 67600 16184 67900 6 wbs_cyc_i
port 348 nsew signal input
rlabel metal3 s 59600 60144 59900 60200 6 wbs_dat_i[0]
port 349 nsew signal input
rlabel metal3 s 100 49056 400 49112 6 wbs_dat_i[10]
port 350 nsew signal input
rlabel metal3 s 100 54096 400 54152 6 wbs_dat_i[11]
port 351 nsew signal input
rlabel metal3 s 100 51744 400 51800 6 wbs_dat_i[12]
port 352 nsew signal input
rlabel metal2 s 2352 100 2408 400 6 wbs_dat_i[13]
port 353 nsew signal input
rlabel metal3 s 100 13440 400 13496 6 wbs_dat_i[14]
port 354 nsew signal input
rlabel metal3 s 59600 37968 59900 38024 6 wbs_dat_i[15]
port 355 nsew signal input
rlabel metal2 s 36960 100 37016 400 6 wbs_dat_i[16]
port 356 nsew signal input
rlabel metal2 s 39648 67600 39704 67900 6 wbs_dat_i[17]
port 357 nsew signal input
rlabel metal2 s 55104 67600 55160 67900 6 wbs_dat_i[18]
port 358 nsew signal input
rlabel metal3 s 100 67872 400 67928 6 wbs_dat_i[19]
port 359 nsew signal input
rlabel metal2 s 9744 100 9800 400 6 wbs_dat_i[1]
port 360 nsew signal input
rlabel metal3 s 100 29904 400 29960 6 wbs_dat_i[20]
port 361 nsew signal input
rlabel metal2 s 56784 67600 56840 67900 6 wbs_dat_i[21]
port 362 nsew signal input
rlabel metal3 s 100 37968 400 38024 6 wbs_dat_i[22]
port 363 nsew signal input
rlabel metal3 s 59600 54432 59900 54488 6 wbs_dat_i[23]
port 364 nsew signal input
rlabel metal3 s 59600 24864 59900 24920 6 wbs_dat_i[24]
port 365 nsew signal input
rlabel metal2 s 44352 100 44408 400 6 wbs_dat_i[25]
port 366 nsew signal input
rlabel metal2 s 49392 67600 49448 67900 6 wbs_dat_i[26]
port 367 nsew signal input
rlabel metal2 s 11088 67600 11144 67900 6 wbs_dat_i[27]
port 368 nsew signal input
rlabel metal2 s 20160 100 20216 400 6 wbs_dat_i[28]
port 369 nsew signal input
rlabel metal3 s 59600 42672 59900 42728 6 wbs_dat_i[29]
port 370 nsew signal input
rlabel metal2 s 52416 100 52472 400 6 wbs_dat_i[2]
port 371 nsew signal input
rlabel metal3 s 59600 22848 59900 22904 6 wbs_dat_i[30]
port 372 nsew signal input
rlabel metal3 s 100 33936 400 33992 6 wbs_dat_i[31]
port 373 nsew signal input
rlabel metal3 s 59600 6384 59900 6440 6 wbs_dat_i[3]
port 374 nsew signal input
rlabel metal2 s 10416 100 10472 400 6 wbs_dat_i[4]
port 375 nsew signal input
rlabel metal2 s 31920 100 31976 400 6 wbs_dat_i[5]
port 376 nsew signal input
rlabel metal3 s 59600 31584 59900 31640 6 wbs_dat_i[6]
port 377 nsew signal input
rlabel metal2 s 46368 67600 46424 67900 6 wbs_dat_i[7]
port 378 nsew signal input
rlabel metal3 s 59600 61152 59900 61208 6 wbs_dat_i[8]
port 379 nsew signal input
rlabel metal3 s 59600 7728 59900 7784 6 wbs_dat_i[9]
port 380 nsew signal input
rlabel metal3 s 100 12768 400 12824 6 wbs_dat_o[0]
port 381 nsew signal output
rlabel metal3 s 59600 40992 59900 41048 6 wbs_dat_o[10]
port 382 nsew signal output
rlabel metal2 s 1008 100 1064 400 6 wbs_dat_o[11]
port 383 nsew signal output
rlabel metal3 s 59600 63168 59900 63224 6 wbs_dat_o[12]
port 384 nsew signal output
rlabel metal2 s 44016 67600 44072 67900 6 wbs_dat_o[13]
port 385 nsew signal output
rlabel metal3 s 59600 11424 59900 11480 6 wbs_dat_o[14]
port 386 nsew signal output
rlabel metal2 s 42000 67600 42056 67900 6 wbs_dat_o[15]
port 387 nsew signal output
rlabel metal3 s 100 17808 400 17864 6 wbs_dat_o[16]
port 388 nsew signal output
rlabel metal3 s 100 20160 400 20216 6 wbs_dat_o[17]
port 389 nsew signal output
rlabel metal2 s 43008 100 43064 400 6 wbs_dat_o[18]
port 390 nsew signal output
rlabel metal2 s 0 100 56 400 6 wbs_dat_o[19]
port 391 nsew signal output
rlabel metal2 s 50400 100 50456 400 6 wbs_dat_o[1]
port 392 nsew signal output
rlabel metal3 s 100 30576 400 30632 6 wbs_dat_o[20]
port 393 nsew signal output
rlabel metal3 s 100 55440 400 55496 6 wbs_dat_o[21]
port 394 nsew signal output
rlabel metal2 s 13776 67600 13832 67900 6 wbs_dat_o[22]
port 395 nsew signal output
rlabel metal3 s 100 20832 400 20888 6 wbs_dat_o[23]
port 396 nsew signal output
rlabel metal2 s 13440 100 13496 400 6 wbs_dat_o[24]
port 397 nsew signal output
rlabel metal2 s 4704 100 4760 400 6 wbs_dat_o[25]
port 398 nsew signal output
rlabel metal2 s 29232 67600 29288 67900 6 wbs_dat_o[26]
port 399 nsew signal output
rlabel metal2 s 14784 67600 14840 67900 6 wbs_dat_o[27]
port 400 nsew signal output
rlabel metal2 s 34944 100 35000 400 6 wbs_dat_o[28]
port 401 nsew signal output
rlabel metal2 s 40320 67600 40376 67900 6 wbs_dat_o[29]
port 402 nsew signal output
rlabel metal3 s 59600 21840 59900 21896 6 wbs_dat_o[2]
port 403 nsew signal output
rlabel metal3 s 100 41664 400 41720 6 wbs_dat_o[30]
port 404 nsew signal output
rlabel metal3 s 59600 53760 59900 53816 6 wbs_dat_o[31]
port 405 nsew signal output
rlabel metal2 s 14112 100 14168 400 6 wbs_dat_o[3]
port 406 nsew signal output
rlabel metal2 s 24528 100 24584 400 6 wbs_dat_o[4]
port 407 nsew signal output
rlabel metal3 s 100 5376 400 5432 6 wbs_dat_o[5]
port 408 nsew signal output
rlabel metal3 s 59600 51408 59900 51464 6 wbs_dat_o[6]
port 409 nsew signal output
rlabel metal2 s 38640 100 38696 400 6 wbs_dat_o[7]
port 410 nsew signal output
rlabel metal2 s 37632 67600 37688 67900 6 wbs_dat_o[8]
port 411 nsew signal output
rlabel metal2 s 37296 67600 37352 67900 6 wbs_dat_o[9]
port 412 nsew signal output
rlabel metal3 s 100 59136 400 59192 6 wbs_sel_i[0]
port 413 nsew signal input
rlabel metal2 s 2688 67600 2744 67900 6 wbs_sel_i[1]
port 414 nsew signal input
rlabel metal2 s 46032 100 46088 400 6 wbs_sel_i[2]
port 415 nsew signal input
rlabel metal3 s 100 14112 400 14168 6 wbs_sel_i[3]
port 416 nsew signal input
rlabel metal3 s 100 52752 400 52808 6 wbs_stb_i
port 417 nsew signal input
rlabel metal3 s 59600 35280 59900 35336 6 wbs_we_i
port 418 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 60000 68000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1740154
string GDS_FILE /home/runner/work/tiny_user_project_xls_popcount/tiny_user_project_xls_popcount/openlane/tiny_user_project/runs/22_12_05_08_30/results/signoff/tiny_user_project.magic.gds
string GDS_START 105924
<< end >>

